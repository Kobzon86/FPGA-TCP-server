// ethernet_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ethernet_sys (
		input  wire        clk_50_clk,                             //                        clk_50.clk
		input  wire        clk_ref_125_clk,                        //                   clk_ref_125.clk
		output wire        eth_tse_0_mac_mdio_connection_mdc,      // eth_tse_0_mac_mdio_connection.mdc
		input  wire        eth_tse_0_mac_mdio_connection_mdio_in,  //                              .mdio_in
		output wire        eth_tse_0_mac_mdio_connection_mdio_out, //                              .mdio_out
		output wire        eth_tse_0_mac_mdio_connection_mdio_oen, //                              .mdio_oen
		output wire        lcd_16207_0_external_RS,                //          lcd_16207_0_external.RS
		output wire        lcd_16207_0_external_RW,                //                              .RW
		inout  wire [7:0]  lcd_16207_0_external_data,              //                              .data
		output wire        lcd_16207_0_external_E,                 //                              .E
		output wire        leds_crs,                               //                          leds.crs
		output wire        leds_link,                              //                              .link
		output wire        leds_panel_link,                        //                              .panel_link
		output wire        leds_col,                               //                              .col
		output wire        leds_an,                                //                              .an
		output wire        leds_char_err,                          //                              .char_err
		output wire        leds_disp_err,                          //                              .disp_err
		input  wire        mac_misc_ff_tx_crc_fwd,                 //                      mac_misc.ff_tx_crc_fwd
		output wire        mac_misc_ff_tx_septy,                   //                              .ff_tx_septy
		output wire        mac_misc_tx_ff_uflow,                   //                              .tx_ff_uflow
		output wire        mac_misc_ff_tx_a_full,                  //                              .ff_tx_a_full
		output wire        mac_misc_ff_tx_a_empty,                 //                              .ff_tx_a_empty
		output wire [17:0] mac_misc_rx_err_stat,                   //                              .rx_err_stat
		output wire [3:0]  mac_misc_rx_frm_type,                   //                              .rx_frm_type
		output wire        mac_misc_ff_rx_dsav,                    //                              .ff_rx_dsav
		output wire        mac_misc_ff_rx_a_full,                  //                              .ff_rx_a_full
		output wire        mac_misc_ff_rx_a_empty,                 //                              .ff_rx_a_empty
		input  wire [7:0]  pio_0_external_connection_export,       //     pio_0_external_connection.export
		output wire [2:0]  pio_1_external_connection_export,       //     pio_1_external_connection.export
		input  wire        reset_reset_n,                          //                         reset.reset_n
		input  wire        reset_0_reset_n,                        //                       reset_0.reset_n
		output wire        serdes_txp,                             //                        serdes.txp
		input  wire        serdes_rxp,                             //                              .rxp
		output wire        serdes_control_rx_recovclkout,          //                serdes_control.rx_recovclkout
		input  wire        serdes_control_reconfig_clk,            //                              .reconfig_clk
		input  wire [3:0]  serdes_control_reconfig_togxb,          //                              .reconfig_togxb
		output wire [4:0]  serdes_control_reconfig_fromgxb,        //                              .reconfig_fromgxb
		input  wire        serdes_control_reconfig_busy,           //                              .reconfig_busy
		output wire        sram_clk_clk,                           //                      sram_clk.clk
		inout  wire [15:0] sram_cntrlr_0_conduit_end_dq,           //     sram_cntrlr_0_conduit_end.dq
		output wire [20:0] sram_cntrlr_0_conduit_end_addr,         //                              .addr
		output wire        sram_cntrlr_0_conduit_end_sram_bwan,    //                              .sram_bwan
		output wire        sram_cntrlr_0_conduit_end_sram_bwbn,    //                              .sram_bwbn
		output wire        sram_cntrlr_0_conduit_end_sram_cen,     //                              .sram_cen
		output wire        sram_cntrlr_0_conduit_end_sram_oen,     //                              .sram_oen
		output wire        sram_cntrlr_0_conduit_end_sram_wen      //                              .sram_wen
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [21:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [21:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sram_cntrlr_0_avalon_slave_readdata;       // sram_cntrlr_0:avalon_slave_readdata -> mm_interconnect_0:sram_cntrlr_0_avalon_slave_readdata
	wire         mm_interconnect_0_sram_cntrlr_0_avalon_slave_waitrequest;    // sram_cntrlr_0:avalon_slave_waitrequest -> mm_interconnect_0:sram_cntrlr_0_avalon_slave_waitrequest
	wire  [18:0] mm_interconnect_0_sram_cntrlr_0_avalon_slave_address;        // mm_interconnect_0:sram_cntrlr_0_avalon_slave_address -> sram_cntrlr_0:avalon_slave_address
	wire         mm_interconnect_0_sram_cntrlr_0_avalon_slave_read;           // mm_interconnect_0:sram_cntrlr_0_avalon_slave_read -> sram_cntrlr_0:avalon_slave_read
	wire   [3:0] mm_interconnect_0_sram_cntrlr_0_avalon_slave_byteenable;     // mm_interconnect_0:sram_cntrlr_0_avalon_slave_byteenable -> sram_cntrlr_0:avalon_slave_byteenable
	wire         mm_interconnect_0_sram_cntrlr_0_avalon_slave_readdatavalid;  // sram_cntrlr_0:avalon_slave_readdatavalid -> mm_interconnect_0:sram_cntrlr_0_avalon_slave_readdatavalid
	wire         mm_interconnect_0_sram_cntrlr_0_avalon_slave_write;          // mm_interconnect_0:sram_cntrlr_0_avalon_slave_write -> sram_cntrlr_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_sram_cntrlr_0_avalon_slave_writedata;      // mm_interconnect_0:sram_cntrlr_0_avalon_slave_writedata -> sram_cntrlr_0:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_eth_tse_0_control_port_readdata;           // eth_tse_0:reg_data_out -> mm_interconnect_0:eth_tse_0_control_port_readdata
	wire         mm_interconnect_0_eth_tse_0_control_port_waitrequest;        // eth_tse_0:reg_busy -> mm_interconnect_0:eth_tse_0_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_eth_tse_0_control_port_address;            // mm_interconnect_0:eth_tse_0_control_port_address -> eth_tse_0:reg_addr
	wire         mm_interconnect_0_eth_tse_0_control_port_read;               // mm_interconnect_0:eth_tse_0_control_port_read -> eth_tse_0:reg_rd
	wire         mm_interconnect_0_eth_tse_0_control_port_write;              // mm_interconnect_0:eth_tse_0_control_port_write -> eth_tse_0:reg_wr
	wire  [31:0] mm_interconnect_0_eth_tse_0_control_port_writedata;          // mm_interconnect_0:eth_tse_0_control_port_writedata -> eth_tse_0:reg_data_in
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_readdata;        // lcd_16207_0:readdata -> mm_interconnect_0:lcd_16207_0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_16207_0_control_slave_address;         // mm_interconnect_0:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	wire         mm_interconnect_0_lcd_16207_0_control_slave_read;            // mm_interconnect_0:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	wire         mm_interconnect_0_lcd_16207_0_control_slave_begintransfer;   // mm_interconnect_0:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	wire         mm_interconnect_0_lcd_16207_0_control_slave_write;           // mm_interconnect_0:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_writedata;       // mm_interconnect_0:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	wire         mm_interconnect_0_sgdma_0_csr_chipselect;                    // mm_interconnect_0:sgdma_0_csr_chipselect -> sgdma_0:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_0_csr_readdata;                      // sgdma_0:csr_readdata -> mm_interconnect_0:sgdma_0_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_0_csr_address;                       // mm_interconnect_0:sgdma_0_csr_address -> sgdma_0:csr_address
	wire         mm_interconnect_0_sgdma_0_csr_read;                          // mm_interconnect_0:sgdma_0_csr_read -> sgdma_0:csr_read
	wire         mm_interconnect_0_sgdma_0_csr_write;                         // mm_interconnect_0:sgdma_0_csr_write -> sgdma_0:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_0_csr_writedata;                     // mm_interconnect_0:sgdma_0_csr_writedata -> sgdma_0:csr_writedata
	wire         mm_interconnect_0_sgdma_1_csr_chipselect;                    // mm_interconnect_0:sgdma_1_csr_chipselect -> sgdma_1:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_1_csr_readdata;                      // sgdma_1:csr_readdata -> mm_interconnect_0:sgdma_1_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_1_csr_address;                       // mm_interconnect_0:sgdma_1_csr_address -> sgdma_1:csr_address
	wire         mm_interconnect_0_sgdma_1_csr_read;                          // mm_interconnect_0:sgdma_1_csr_read -> sgdma_1:csr_read
	wire         mm_interconnect_0_sgdma_1_csr_write;                         // mm_interconnect_0:sgdma_1_csr_write -> sgdma_1:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_1_csr_writedata;                     // mm_interconnect_0:sgdma_1_csr_writedata -> sgdma_1:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                         // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                          // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_pio_1_s1_chipselect;                       // mm_interconnect_0:pio_1_s1_chipselect -> pio_1:chipselect
	wire  [31:0] mm_interconnect_0_pio_1_s1_readdata;                         // pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_1_s1_address;                          // mm_interconnect_0:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_0_pio_1_s1_write;                            // mm_interconnect_0:pio_1_s1_write -> pio_1:write_n
	wire  [31:0] mm_interconnect_0_pio_1_s1_writedata;                        // mm_interconnect_0:pio_1_s1_writedata -> pio_1:writedata
	wire         mm_interconnect_0_descriptor_memory_s2_chipselect;           // mm_interconnect_0:descriptor_memory_s2_chipselect -> descriptor_memory:chipselect2
	wire  [31:0] mm_interconnect_0_descriptor_memory_s2_readdata;             // descriptor_memory:readdata2 -> mm_interconnect_0:descriptor_memory_s2_readdata
	wire   [9:0] mm_interconnect_0_descriptor_memory_s2_address;              // mm_interconnect_0:descriptor_memory_s2_address -> descriptor_memory:address2
	wire   [3:0] mm_interconnect_0_descriptor_memory_s2_byteenable;           // mm_interconnect_0:descriptor_memory_s2_byteenable -> descriptor_memory:byteenable2
	wire         mm_interconnect_0_descriptor_memory_s2_write;                // mm_interconnect_0:descriptor_memory_s2_write -> descriptor_memory:write2
	wire  [31:0] mm_interconnect_0_descriptor_memory_s2_writedata;            // mm_interconnect_0:descriptor_memory_s2_writedata -> descriptor_memory:writedata2
	wire         mm_interconnect_0_descriptor_memory_s2_clken;                // mm_interconnect_0:descriptor_memory_s2_clken -> descriptor_memory:clken2
	wire         mm_interconnect_0_onchip_memory2_0_s2_chipselect;            // mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s2_readdata;              // onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s2_address;               // mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s2_byteenable;            // mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire         mm_interconnect_0_onchip_memory2_0_s2_write;                 // mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s2_writedata;             // mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_0_onchip_memory2_0_s2_clken;                 // mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire  [31:0] sgdma_1_descriptor_read_readdata;                            // mm_interconnect_1:sgdma_1_descriptor_read_readdata -> sgdma_1:descriptor_read_readdata
	wire         sgdma_1_descriptor_read_waitrequest;                         // mm_interconnect_1:sgdma_1_descriptor_read_waitrequest -> sgdma_1:descriptor_read_waitrequest
	wire  [31:0] sgdma_1_descriptor_read_address;                             // sgdma_1:descriptor_read_address -> mm_interconnect_1:sgdma_1_descriptor_read_address
	wire         sgdma_1_descriptor_read_read;                                // sgdma_1:descriptor_read_read -> mm_interconnect_1:sgdma_1_descriptor_read_read
	wire         sgdma_1_descriptor_read_readdatavalid;                       // mm_interconnect_1:sgdma_1_descriptor_read_readdatavalid -> sgdma_1:descriptor_read_readdatavalid
	wire  [31:0] sgdma_0_descriptor_read_readdata;                            // mm_interconnect_1:sgdma_0_descriptor_read_readdata -> sgdma_0:descriptor_read_readdata
	wire         sgdma_0_descriptor_read_waitrequest;                         // mm_interconnect_1:sgdma_0_descriptor_read_waitrequest -> sgdma_0:descriptor_read_waitrequest
	wire  [31:0] sgdma_0_descriptor_read_address;                             // sgdma_0:descriptor_read_address -> mm_interconnect_1:sgdma_0_descriptor_read_address
	wire         sgdma_0_descriptor_read_read;                                // sgdma_0:descriptor_read_read -> mm_interconnect_1:sgdma_0_descriptor_read_read
	wire         sgdma_0_descriptor_read_readdatavalid;                       // mm_interconnect_1:sgdma_0_descriptor_read_readdatavalid -> sgdma_0:descriptor_read_readdatavalid
	wire         sgdma_1_descriptor_write_waitrequest;                        // mm_interconnect_1:sgdma_1_descriptor_write_waitrequest -> sgdma_1:descriptor_write_waitrequest
	wire  [31:0] sgdma_1_descriptor_write_address;                            // sgdma_1:descriptor_write_address -> mm_interconnect_1:sgdma_1_descriptor_write_address
	wire         sgdma_1_descriptor_write_write;                              // sgdma_1:descriptor_write_write -> mm_interconnect_1:sgdma_1_descriptor_write_write
	wire  [31:0] sgdma_1_descriptor_write_writedata;                          // sgdma_1:descriptor_write_writedata -> mm_interconnect_1:sgdma_1_descriptor_write_writedata
	wire         sgdma_0_descriptor_write_waitrequest;                        // mm_interconnect_1:sgdma_0_descriptor_write_waitrequest -> sgdma_0:descriptor_write_waitrequest
	wire  [31:0] sgdma_0_descriptor_write_address;                            // sgdma_0:descriptor_write_address -> mm_interconnect_1:sgdma_0_descriptor_write_address
	wire         sgdma_0_descriptor_write_write;                              // sgdma_0:descriptor_write_write -> mm_interconnect_1:sgdma_0_descriptor_write_write
	wire  [31:0] sgdma_0_descriptor_write_writedata;                          // sgdma_0:descriptor_write_writedata -> mm_interconnect_1:sgdma_0_descriptor_write_writedata
	wire         mm_interconnect_1_descriptor_memory_s1_chipselect;           // mm_interconnect_1:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_readdata;             // descriptor_memory:readdata -> mm_interconnect_1:descriptor_memory_s1_readdata
	wire   [9:0] mm_interconnect_1_descriptor_memory_s1_address;              // mm_interconnect_1:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_1_descriptor_memory_s1_byteenable;           // mm_interconnect_1:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_1_descriptor_memory_s1_write;                // mm_interconnect_1:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_writedata;            // mm_interconnect_1:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_1_descriptor_memory_s1_clken;                // mm_interconnect_1:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire  [31:0] sgdma_0_m_read_readdata;                                     // mm_interconnect_2:sgdma_0_m_read_readdata -> sgdma_0:m_read_readdata
	wire         sgdma_0_m_read_waitrequest;                                  // mm_interconnect_2:sgdma_0_m_read_waitrequest -> sgdma_0:m_read_waitrequest
	wire  [31:0] sgdma_0_m_read_address;                                      // sgdma_0:m_read_address -> mm_interconnect_2:sgdma_0_m_read_address
	wire         sgdma_0_m_read_read;                                         // sgdma_0:m_read_read -> mm_interconnect_2:sgdma_0_m_read_read
	wire         sgdma_0_m_read_readdatavalid;                                // mm_interconnect_2:sgdma_0_m_read_readdatavalid -> sgdma_0:m_read_readdatavalid
	wire         sgdma_1_m_write_waitrequest;                                 // mm_interconnect_2:sgdma_1_m_write_waitrequest -> sgdma_1:m_write_waitrequest
	wire  [31:0] sgdma_1_m_write_address;                                     // sgdma_1:m_write_address -> mm_interconnect_2:sgdma_1_m_write_address
	wire   [3:0] sgdma_1_m_write_byteenable;                                  // sgdma_1:m_write_byteenable -> mm_interconnect_2:sgdma_1_m_write_byteenable
	wire         sgdma_1_m_write_write;                                       // sgdma_1:m_write_write -> mm_interconnect_2:sgdma_1_m_write_write
	wire  [31:0] sgdma_1_m_write_writedata;                                   // sgdma_1:m_write_writedata -> mm_interconnect_2:sgdma_1_m_write_writedata
	wire         mm_interconnect_2_onchip_memory2_0_s1_chipselect;            // mm_interconnect_2:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_2_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_2:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_2_onchip_memory2_0_s1_address;               // mm_interconnect_2:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_2_onchip_memory2_0_s1_byteenable;            // mm_interconnect_2:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_2_onchip_memory2_0_s1_write;                 // mm_interconnect_2:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_2_onchip_memory2_0_s1_writedata;             // mm_interconnect_2:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_2_onchip_memory2_0_s1_clken;                 // mm_interconnect_2:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                    // sgdma_1:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // sgdma_0:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         sgdma_0_out_valid;                                           // sgdma_0:out_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] sgdma_0_out_data;                                            // sgdma_0:out_data -> avalon_st_adapter:in_0_data
	wire         sgdma_0_out_ready;                                           // avalon_st_adapter:in_0_ready -> sgdma_0:out_ready
	wire         sgdma_0_out_startofpacket;                                   // sgdma_0:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         sgdma_0_out_endofpacket;                                     // sgdma_0:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire   [1:0] sgdma_0_out_empty;                                           // sgdma_0:out_empty -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                               // avalon_st_adapter:out_0_valid -> eth_tse_0:ff_tx_wren
	wire  [31:0] avalon_st_adapter_out_0_data;                                // avalon_st_adapter:out_0_data -> eth_tse_0:ff_tx_data
	wire         avalon_st_adapter_out_0_ready;                               // eth_tse_0:ff_tx_rdy -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                       // avalon_st_adapter:out_0_startofpacket -> eth_tse_0:ff_tx_sop
	wire         avalon_st_adapter_out_0_endofpacket;                         // avalon_st_adapter:out_0_endofpacket -> eth_tse_0:ff_tx_eop
	wire   [0:0] avalon_st_adapter_out_0_error;                               // avalon_st_adapter:out_0_error -> eth_tse_0:ff_tx_err
	wire   [1:0] avalon_st_adapter_out_0_empty;                               // avalon_st_adapter:out_0_empty -> eth_tse_0:ff_tx_mod
	wire         eth_tse_0_receive_valid;                                     // eth_tse_0:ff_rx_dval -> avalon_st_adapter_001:in_0_valid
	wire  [31:0] eth_tse_0_receive_data;                                      // eth_tse_0:ff_rx_data -> avalon_st_adapter_001:in_0_data
	wire         eth_tse_0_receive_ready;                                     // avalon_st_adapter_001:in_0_ready -> eth_tse_0:ff_rx_rdy
	wire         eth_tse_0_receive_startofpacket;                             // eth_tse_0:ff_rx_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire         eth_tse_0_receive_endofpacket;                               // eth_tse_0:ff_rx_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire   [5:0] eth_tse_0_receive_error;                                     // eth_tse_0:rx_err -> avalon_st_adapter_001:in_0_error
	wire   [1:0] eth_tse_0_receive_empty;                                     // eth_tse_0:ff_rx_mod -> avalon_st_adapter_001:in_0_empty
	wire         avalon_st_adapter_001_out_0_valid;                           // avalon_st_adapter_001:out_0_valid -> sgdma_1:in_valid
	wire  [31:0] avalon_st_adapter_001_out_0_data;                            // avalon_st_adapter_001:out_0_data -> sgdma_1:in_data
	wire         avalon_st_adapter_001_out_0_ready;                           // sgdma_1:in_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;                   // avalon_st_adapter_001:out_0_startofpacket -> sgdma_1:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                     // avalon_st_adapter_001:out_0_endofpacket -> sgdma_1:in_endofpacket
	wire   [1:0] avalon_st_adapter_001_out_0_empty;                           // avalon_st_adapter_001:out_0_empty -> sgdma_1:in_empty
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> altpll_0:reset
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, descriptor_memory:reset, eth_tse_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, lcd_16207_0:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sgdma_1_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sgdma_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, pio_0:reset_n, pio_1:reset_n, rst_translator:in_reset, sgdma_0:system_reset_n, sgdma_1:system_reset_n, sram_cntrlr_0:rst_n, timer_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [descriptor_memory:reset_req, nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	ethernet_sys_altpll_0 altpll_0 (
		.clk                (clk_50_clk),                     //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (sram_clk_clk),                   //                    c0.clk
		.locked             (),                               //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.areset             (1'b0),                           //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (4'b0000),                        //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	ethernet_sys_descriptor_memory descriptor_memory (
		.address     (mm_interconnect_1_descriptor_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_descriptor_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_descriptor_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_descriptor_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_1_descriptor_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_descriptor_memory_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_descriptor_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_descriptor_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_descriptor_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_descriptor_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_descriptor_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_descriptor_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_descriptor_memory_s2_byteenable), //       .byteenable
		.clk         (sram_clk_clk),                                      //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),            //       .reset_req
		.freeze      (1'b0)                                               // (terminated)
	);

	ethernet_sys_eth_tse_0 eth_tse_0 (
		.clk              (sram_clk_clk),                                         // control_port_clock_connection.clk
		.reset            (rst_controller_001_reset_out_reset),                   //              reset_connection.reset
		.reg_data_out     (mm_interconnect_0_eth_tse_0_control_port_readdata),    //                  control_port.readdata
		.reg_rd           (mm_interconnect_0_eth_tse_0_control_port_read),        //                              .read
		.reg_data_in      (mm_interconnect_0_eth_tse_0_control_port_writedata),   //                              .writedata
		.reg_wr           (mm_interconnect_0_eth_tse_0_control_port_write),       //                              .write
		.reg_busy         (mm_interconnect_0_eth_tse_0_control_port_waitrequest), //                              .waitrequest
		.reg_addr         (mm_interconnect_0_eth_tse_0_control_port_address),     //                              .address
		.ff_rx_clk        (sram_clk_clk),                                         //      receive_clock_connection.clk
		.ff_tx_clk        (sram_clk_clk),                                         //     transmit_clock_connection.clk
		.ff_rx_data       (eth_tse_0_receive_data),                               //                       receive.data
		.ff_rx_eop        (eth_tse_0_receive_endofpacket),                        //                              .endofpacket
		.rx_err           (eth_tse_0_receive_error),                              //                              .error
		.ff_rx_mod        (eth_tse_0_receive_empty),                              //                              .empty
		.ff_rx_rdy        (eth_tse_0_receive_ready),                              //                              .ready
		.ff_rx_sop        (eth_tse_0_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval       (eth_tse_0_receive_valid),                              //                              .valid
		.ff_tx_data       (avalon_st_adapter_out_0_data),                         //                      transmit.data
		.ff_tx_eop        (avalon_st_adapter_out_0_endofpacket),                  //                              .endofpacket
		.ff_tx_err        (avalon_st_adapter_out_0_error),                        //                              .error
		.ff_tx_mod        (avalon_st_adapter_out_0_empty),                        //                              .empty
		.ff_tx_rdy        (avalon_st_adapter_out_0_ready),                        //                              .ready
		.ff_tx_sop        (avalon_st_adapter_out_0_startofpacket),                //                              .startofpacket
		.ff_tx_wren       (avalon_st_adapter_out_0_valid),                        //                              .valid
		.mdc              (eth_tse_0_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in          (eth_tse_0_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out         (eth_tse_0_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen         (eth_tse_0_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.ff_tx_crc_fwd    (mac_misc_ff_tx_crc_fwd),                               //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy      (mac_misc_ff_tx_septy),                                 //                              .ff_tx_septy
		.tx_ff_uflow      (mac_misc_tx_ff_uflow),                                 //                              .tx_ff_uflow
		.ff_tx_a_full     (mac_misc_ff_tx_a_full),                                //                              .ff_tx_a_full
		.ff_tx_a_empty    (mac_misc_ff_tx_a_empty),                               //                              .ff_tx_a_empty
		.rx_err_stat      (mac_misc_rx_err_stat),                                 //                              .rx_err_stat
		.rx_frm_type      (mac_misc_rx_frm_type),                                 //                              .rx_frm_type
		.ff_rx_dsav       (mac_misc_ff_rx_dsav),                                  //                              .ff_rx_dsav
		.ff_rx_a_full     (mac_misc_ff_rx_a_full),                                //                              .ff_rx_a_full
		.ff_rx_a_empty    (mac_misc_ff_rx_a_empty),                               //                              .ff_rx_a_empty
		.ref_clk          (clk_ref_125_clk),                                      //  pcs_ref_clk_clock_connection.clk
		.gxb_cal_blk_clk  (sram_clk_clk),                                         //                   cal_blk_clk.clk
		.led_crs          (leds_crs),                                             //         status_led_connection.crs
		.led_link         (leds_link),                                            //                              .link
		.led_panel_link   (leds_panel_link),                                      //                              .panel_link
		.led_col          (leds_col),                                             //                              .col
		.led_an           (leds_an),                                              //                              .an
		.led_char_err     (leds_char_err),                                        //                              .char_err
		.led_disp_err     (leds_disp_err),                                        //                              .disp_err
		.rx_recovclkout   (serdes_control_rx_recovclkout),                        //     serdes_control_connection.rx_recovclkout
		.reconfig_clk     (serdes_control_reconfig_clk),                          //                              .reconfig_clk
		.reconfig_togxb   (serdes_control_reconfig_togxb),                        //                              .reconfig_togxb
		.reconfig_fromgxb (serdes_control_reconfig_fromgxb),                      //                              .reconfig_fromgxb
		.reconfig_busy    (serdes_control_reconfig_busy),                         //                              .reconfig_busy
		.txp              (serdes_txp),                                           //             serial_connection.txp
		.rxp              (serdes_rxp)                                            //                              .rxp
	);

	ethernet_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (sram_clk_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	ethernet_sys_lcd_16207_0 lcd_16207_0 (
		.reset_n       (~rst_controller_001_reset_out_reset),                       //         reset.reset_n
		.clk           (sram_clk_clk),                                              //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_16207_0_external_RS),                                   //      external.export
		.LCD_RW        (lcd_16207_0_external_RW),                                   //              .export
		.LCD_data      (lcd_16207_0_external_data),                                 //              .export
		.LCD_E         (lcd_16207_0_external_E)                                     //              .export
	);

	ethernet_sys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sram_clk_clk),                                               //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	ethernet_sys_onchip_memory2_0 onchip_memory2_0 (
		.address     (mm_interconnect_2_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_2_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_onchip_memory2_0_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk         (sram_clk_clk),                                     //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	ethernet_sys_pio_0 pio_0 (
		.clk      (sram_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_pio_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_0_s1_readdata), //                    .readdata
		.in_port  (pio_0_external_connection_export)     // external_connection.export
	);

	ethernet_sys_pio_1 pio_1 (
		.clk        (sram_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_pio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_1_s1_readdata),   //                    .readdata
		.out_port   (pio_1_external_connection_export)       // external_connection.export
	);

	ethernet_sys_sgdma_0 sgdma_0 (
		.clk                           (sram_clk_clk),                             //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),      //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_0_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_0_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_0_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_0_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_0_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_0_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_0_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_0_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_0_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_0_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_0_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_0_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_0_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_0_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_0_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                 //          csr_irq.irq
		.m_read_readdata               (sgdma_0_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_0_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_0_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_0_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_0_m_read_read),                      //                 .read
		.out_data                      (sgdma_0_out_data),                         //              out.data
		.out_valid                     (sgdma_0_out_valid),                        //                 .valid
		.out_ready                     (sgdma_0_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_0_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_0_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_0_out_empty)                         //                 .empty
	);

	ethernet_sys_sgdma_1 sgdma_1 (
		.clk                           (sram_clk_clk),                              //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_1_csr_chipselect),  //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_1_csr_address),     //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_1_csr_read),        //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_1_csr_write),       //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_1_csr_writedata),   //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_1_csr_readdata),    //                 .readdata
		.descriptor_read_readdata      (sgdma_1_descriptor_read_readdata),          //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_1_descriptor_read_readdatavalid),     //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_1_descriptor_read_waitrequest),       //                 .waitrequest
		.descriptor_read_address       (sgdma_1_descriptor_read_address),           //                 .address
		.descriptor_read_read          (sgdma_1_descriptor_read_read),              //                 .read
		.descriptor_write_waitrequest  (sgdma_1_descriptor_write_waitrequest),      // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_1_descriptor_write_address),          //                 .address
		.descriptor_write_write        (sgdma_1_descriptor_write_write),            //                 .write
		.descriptor_write_writedata    (sgdma_1_descriptor_write_writedata),        //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_001_out_0_startofpacket), //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_001_out_0_endofpacket),   //                 .endofpacket
		.in_data                       (avalon_st_adapter_001_out_0_data),          //                 .data
		.in_valid                      (avalon_st_adapter_001_out_0_valid),         //                 .valid
		.in_ready                      (avalon_st_adapter_001_out_0_ready),         //                 .ready
		.in_empty                      (avalon_st_adapter_001_out_0_empty),         //                 .empty
		.m_write_waitrequest           (sgdma_1_m_write_waitrequest),               //          m_write.waitrequest
		.m_write_address               (sgdma_1_m_write_address),                   //                 .address
		.m_write_write                 (sgdma_1_m_write_write),                     //                 .write
		.m_write_writedata             (sgdma_1_m_write_writedata),                 //                 .writedata
		.m_write_byteenable            (sgdma_1_m_write_byteenable)                 //                 .byteenable
	);

	sram_cntrlr sram_cntrlr_0 (
		.clk                        (sram_clk_clk),                                               //        clock.clk
		.avalon_slave_address       (mm_interconnect_0_sram_cntrlr_0_avalon_slave_address),       // avalon_slave.address
		.avalon_slave_read          (mm_interconnect_0_sram_cntrlr_0_avalon_slave_read),          //             .read
		.avalon_slave_readdata      (mm_interconnect_0_sram_cntrlr_0_avalon_slave_readdata),      //             .readdata
		.avalon_slave_readdatavalid (mm_interconnect_0_sram_cntrlr_0_avalon_slave_readdatavalid), //             .readdatavalid
		.avalon_slave_write         (mm_interconnect_0_sram_cntrlr_0_avalon_slave_write),         //             .write
		.avalon_slave_writedata     (mm_interconnect_0_sram_cntrlr_0_avalon_slave_writedata),     //             .writedata
		.avalon_slave_waitrequest   (mm_interconnect_0_sram_cntrlr_0_avalon_slave_waitrequest),   //             .waitrequest
		.avalon_slave_byteenable    (mm_interconnect_0_sram_cntrlr_0_avalon_slave_byteenable),    //             .byteenable
		.dq                         (sram_cntrlr_0_conduit_end_dq),                               //  conduit_end.dq
		.addr                       (sram_cntrlr_0_conduit_end_addr),                             //             .addr
		.sram_bwan                  (sram_cntrlr_0_conduit_end_sram_bwan),                        //             .sram_bwan
		.sram_bwbn                  (sram_cntrlr_0_conduit_end_sram_bwbn),                        //             .sram_bwbn
		.sram_cen                   (sram_cntrlr_0_conduit_end_sram_cen),                         //             .sram_cen
		.sram_oen                   (sram_cntrlr_0_conduit_end_sram_oen),                         //             .sram_oen
		.sram_wen                   (sram_cntrlr_0_conduit_end_sram_wen),                         //             .sram_wen
		.rst_n                      (~rst_controller_001_reset_out_reset)                         //   reset_sink.reset_n
	);

	ethernet_sys_timer_0 timer_0 (
		.clk        (sram_clk_clk),                            //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	ethernet_sys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                (sram_clk_clk),                                                //                              altpll_0_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.descriptor_memory_s2_address                   (mm_interconnect_0_descriptor_memory_s2_address),              //                     descriptor_memory_s2.address
		.descriptor_memory_s2_write                     (mm_interconnect_0_descriptor_memory_s2_write),                //                                         .write
		.descriptor_memory_s2_readdata                  (mm_interconnect_0_descriptor_memory_s2_readdata),             //                                         .readdata
		.descriptor_memory_s2_writedata                 (mm_interconnect_0_descriptor_memory_s2_writedata),            //                                         .writedata
		.descriptor_memory_s2_byteenable                (mm_interconnect_0_descriptor_memory_s2_byteenable),           //                                         .byteenable
		.descriptor_memory_s2_chipselect                (mm_interconnect_0_descriptor_memory_s2_chipselect),           //                                         .chipselect
		.descriptor_memory_s2_clken                     (mm_interconnect_0_descriptor_memory_s2_clken),                //                                         .clken
		.eth_tse_0_control_port_address                 (mm_interconnect_0_eth_tse_0_control_port_address),            //                   eth_tse_0_control_port.address
		.eth_tse_0_control_port_write                   (mm_interconnect_0_eth_tse_0_control_port_write),              //                                         .write
		.eth_tse_0_control_port_read                    (mm_interconnect_0_eth_tse_0_control_port_read),               //                                         .read
		.eth_tse_0_control_port_readdata                (mm_interconnect_0_eth_tse_0_control_port_readdata),           //                                         .readdata
		.eth_tse_0_control_port_writedata               (mm_interconnect_0_eth_tse_0_control_port_writedata),          //                                         .writedata
		.eth_tse_0_control_port_waitrequest             (mm_interconnect_0_eth_tse_0_control_port_waitrequest),        //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.lcd_16207_0_control_slave_address              (mm_interconnect_0_lcd_16207_0_control_slave_address),         //                lcd_16207_0_control_slave.address
		.lcd_16207_0_control_slave_write                (mm_interconnect_0_lcd_16207_0_control_slave_write),           //                                         .write
		.lcd_16207_0_control_slave_read                 (mm_interconnect_0_lcd_16207_0_control_slave_read),            //                                         .read
		.lcd_16207_0_control_slave_readdata             (mm_interconnect_0_lcd_16207_0_control_slave_readdata),        //                                         .readdata
		.lcd_16207_0_control_slave_writedata            (mm_interconnect_0_lcd_16207_0_control_slave_writedata),       //                                         .writedata
		.lcd_16207_0_control_slave_begintransfer        (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer),   //                                         .begintransfer
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s2_address                    (mm_interconnect_0_onchip_memory2_0_s2_address),               //                      onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                      (mm_interconnect_0_onchip_memory2_0_s2_write),                 //                                         .write
		.onchip_memory2_0_s2_readdata                   (mm_interconnect_0_onchip_memory2_0_s2_readdata),              //                                         .readdata
		.onchip_memory2_0_s2_writedata                  (mm_interconnect_0_onchip_memory2_0_s2_writedata),             //                                         .writedata
		.onchip_memory2_0_s2_byteenable                 (mm_interconnect_0_onchip_memory2_0_s2_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s2_chipselect                 (mm_interconnect_0_onchip_memory2_0_s2_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s2_clken                      (mm_interconnect_0_onchip_memory2_0_s2_clken),                 //                                         .clken
		.pio_0_s1_address                               (mm_interconnect_0_pio_0_s1_address),                          //                                 pio_0_s1.address
		.pio_0_s1_readdata                              (mm_interconnect_0_pio_0_s1_readdata),                         //                                         .readdata
		.pio_1_s1_address                               (mm_interconnect_0_pio_1_s1_address),                          //                                 pio_1_s1.address
		.pio_1_s1_write                                 (mm_interconnect_0_pio_1_s1_write),                            //                                         .write
		.pio_1_s1_readdata                              (mm_interconnect_0_pio_1_s1_readdata),                         //                                         .readdata
		.pio_1_s1_writedata                             (mm_interconnect_0_pio_1_s1_writedata),                        //                                         .writedata
		.pio_1_s1_chipselect                            (mm_interconnect_0_pio_1_s1_chipselect),                       //                                         .chipselect
		.sgdma_0_csr_address                            (mm_interconnect_0_sgdma_0_csr_address),                       //                              sgdma_0_csr.address
		.sgdma_0_csr_write                              (mm_interconnect_0_sgdma_0_csr_write),                         //                                         .write
		.sgdma_0_csr_read                               (mm_interconnect_0_sgdma_0_csr_read),                          //                                         .read
		.sgdma_0_csr_readdata                           (mm_interconnect_0_sgdma_0_csr_readdata),                      //                                         .readdata
		.sgdma_0_csr_writedata                          (mm_interconnect_0_sgdma_0_csr_writedata),                     //                                         .writedata
		.sgdma_0_csr_chipselect                         (mm_interconnect_0_sgdma_0_csr_chipselect),                    //                                         .chipselect
		.sgdma_1_csr_address                            (mm_interconnect_0_sgdma_1_csr_address),                       //                              sgdma_1_csr.address
		.sgdma_1_csr_write                              (mm_interconnect_0_sgdma_1_csr_write),                         //                                         .write
		.sgdma_1_csr_read                               (mm_interconnect_0_sgdma_1_csr_read),                          //                                         .read
		.sgdma_1_csr_readdata                           (mm_interconnect_0_sgdma_1_csr_readdata),                      //                                         .readdata
		.sgdma_1_csr_writedata                          (mm_interconnect_0_sgdma_1_csr_writedata),                     //                                         .writedata
		.sgdma_1_csr_chipselect                         (mm_interconnect_0_sgdma_1_csr_chipselect),                    //                                         .chipselect
		.sram_cntrlr_0_avalon_slave_address             (mm_interconnect_0_sram_cntrlr_0_avalon_slave_address),        //               sram_cntrlr_0_avalon_slave.address
		.sram_cntrlr_0_avalon_slave_write               (mm_interconnect_0_sram_cntrlr_0_avalon_slave_write),          //                                         .write
		.sram_cntrlr_0_avalon_slave_read                (mm_interconnect_0_sram_cntrlr_0_avalon_slave_read),           //                                         .read
		.sram_cntrlr_0_avalon_slave_readdata            (mm_interconnect_0_sram_cntrlr_0_avalon_slave_readdata),       //                                         .readdata
		.sram_cntrlr_0_avalon_slave_writedata           (mm_interconnect_0_sram_cntrlr_0_avalon_slave_writedata),      //                                         .writedata
		.sram_cntrlr_0_avalon_slave_byteenable          (mm_interconnect_0_sram_cntrlr_0_avalon_slave_byteenable),     //                                         .byteenable
		.sram_cntrlr_0_avalon_slave_readdatavalid       (mm_interconnect_0_sram_cntrlr_0_avalon_slave_readdatavalid),  //                                         .readdatavalid
		.sram_cntrlr_0_avalon_slave_waitrequest         (mm_interconnect_0_sram_cntrlr_0_avalon_slave_waitrequest),    //                                         .waitrequest
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                      //                                         .chipselect
	);

	ethernet_sys_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c0_clk                           (sram_clk_clk),                                      //                         altpll_0_c0.clk
		.sgdma_1_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // sgdma_1_reset_reset_bridge_in_reset.reset
		.sgdma_0_descriptor_read_address           (sgdma_0_descriptor_read_address),                   //             sgdma_0_descriptor_read.address
		.sgdma_0_descriptor_read_waitrequest       (sgdma_0_descriptor_read_waitrequest),               //                                    .waitrequest
		.sgdma_0_descriptor_read_read              (sgdma_0_descriptor_read_read),                      //                                    .read
		.sgdma_0_descriptor_read_readdata          (sgdma_0_descriptor_read_readdata),                  //                                    .readdata
		.sgdma_0_descriptor_read_readdatavalid     (sgdma_0_descriptor_read_readdatavalid),             //                                    .readdatavalid
		.sgdma_0_descriptor_write_address          (sgdma_0_descriptor_write_address),                  //            sgdma_0_descriptor_write.address
		.sgdma_0_descriptor_write_waitrequest      (sgdma_0_descriptor_write_waitrequest),              //                                    .waitrequest
		.sgdma_0_descriptor_write_write            (sgdma_0_descriptor_write_write),                    //                                    .write
		.sgdma_0_descriptor_write_writedata        (sgdma_0_descriptor_write_writedata),                //                                    .writedata
		.sgdma_1_descriptor_read_address           (sgdma_1_descriptor_read_address),                   //             sgdma_1_descriptor_read.address
		.sgdma_1_descriptor_read_waitrequest       (sgdma_1_descriptor_read_waitrequest),               //                                    .waitrequest
		.sgdma_1_descriptor_read_read              (sgdma_1_descriptor_read_read),                      //                                    .read
		.sgdma_1_descriptor_read_readdata          (sgdma_1_descriptor_read_readdata),                  //                                    .readdata
		.sgdma_1_descriptor_read_readdatavalid     (sgdma_1_descriptor_read_readdatavalid),             //                                    .readdatavalid
		.sgdma_1_descriptor_write_address          (sgdma_1_descriptor_write_address),                  //            sgdma_1_descriptor_write.address
		.sgdma_1_descriptor_write_waitrequest      (sgdma_1_descriptor_write_waitrequest),              //                                    .waitrequest
		.sgdma_1_descriptor_write_write            (sgdma_1_descriptor_write_write),                    //                                    .write
		.sgdma_1_descriptor_write_writedata        (sgdma_1_descriptor_write_writedata),                //                                    .writedata
		.descriptor_memory_s1_address              (mm_interconnect_1_descriptor_memory_s1_address),    //                descriptor_memory_s1.address
		.descriptor_memory_s1_write                (mm_interconnect_1_descriptor_memory_s1_write),      //                                    .write
		.descriptor_memory_s1_readdata             (mm_interconnect_1_descriptor_memory_s1_readdata),   //                                    .readdata
		.descriptor_memory_s1_writedata            (mm_interconnect_1_descriptor_memory_s1_writedata),  //                                    .writedata
		.descriptor_memory_s1_byteenable           (mm_interconnect_1_descriptor_memory_s1_byteenable), //                                    .byteenable
		.descriptor_memory_s1_chipselect           (mm_interconnect_1_descriptor_memory_s1_chipselect), //                                    .chipselect
		.descriptor_memory_s1_clken                (mm_interconnect_1_descriptor_memory_s1_clken)       //                                    .clken
	);

	ethernet_sys_mm_interconnect_2 mm_interconnect_2 (
		.altpll_0_c0_clk                           (sram_clk_clk),                                     //                         altpll_0_c0.clk
		.sgdma_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),               // sgdma_0_reset_reset_bridge_in_reset.reset
		.sgdma_0_m_read_address                    (sgdma_0_m_read_address),                           //                      sgdma_0_m_read.address
		.sgdma_0_m_read_waitrequest                (sgdma_0_m_read_waitrequest),                       //                                    .waitrequest
		.sgdma_0_m_read_read                       (sgdma_0_m_read_read),                              //                                    .read
		.sgdma_0_m_read_readdata                   (sgdma_0_m_read_readdata),                          //                                    .readdata
		.sgdma_0_m_read_readdatavalid              (sgdma_0_m_read_readdatavalid),                     //                                    .readdatavalid
		.sgdma_1_m_write_address                   (sgdma_1_m_write_address),                          //                     sgdma_1_m_write.address
		.sgdma_1_m_write_waitrequest               (sgdma_1_m_write_waitrequest),                      //                                    .waitrequest
		.sgdma_1_m_write_byteenable                (sgdma_1_m_write_byteenable),                       //                                    .byteenable
		.sgdma_1_m_write_write                     (sgdma_1_m_write_write),                            //                                    .write
		.sgdma_1_m_write_writedata                 (sgdma_1_m_write_writedata),                        //                                    .writedata
		.onchip_memory2_0_s1_address               (mm_interconnect_2_onchip_memory2_0_s1_address),    //                 onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                 (mm_interconnect_2_onchip_memory2_0_s1_write),      //                                    .write
		.onchip_memory2_0_s1_readdata              (mm_interconnect_2_onchip_memory2_0_s1_readdata),   //                                    .readdata
		.onchip_memory2_0_s1_writedata             (mm_interconnect_2_onchip_memory2_0_s1_writedata),  //                                    .writedata
		.onchip_memory2_0_s1_byteenable            (mm_interconnect_2_onchip_memory2_0_s1_byteenable), //                                    .byteenable
		.onchip_memory2_0_s1_chipselect            (mm_interconnect_2_onchip_memory2_0_s1_chipselect), //                                    .chipselect
		.onchip_memory2_0_s1_clken                 (mm_interconnect_2_onchip_memory2_0_s1_clken)       //                                    .clken
	);

	ethernet_sys_irq_mapper irq_mapper (
		.clk           (sram_clk_clk),                       //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	ethernet_sys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sram_clk_clk),                          // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (sgdma_0_out_data),                      //     in_0.data
		.in_0_valid          (sgdma_0_out_valid),                     //         .valid
		.in_0_ready          (sgdma_0_out_ready),                     //         .ready
		.in_0_startofpacket  (sgdma_0_out_startofpacket),             //         .startofpacket
		.in_0_endofpacket    (sgdma_0_out_endofpacket),               //         .endofpacket
		.in_0_empty          (sgdma_0_out_empty),                     //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	ethernet_sys_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (sram_clk_clk),                              // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (eth_tse_0_receive_data),                    //     in_0.data
		.in_0_valid          (eth_tse_0_receive_valid),                   //         .valid
		.in_0_ready          (eth_tse_0_receive_ready),                   //         .ready
		.in_0_startofpacket  (eth_tse_0_receive_startofpacket),           //         .startofpacket
		.in_0_endofpacket    (eth_tse_0_receive_endofpacket),             //         .endofpacket
		.in_0_empty          (eth_tse_0_receive_empty),                   //         .empty
		.in_0_error          (eth_tse_0_receive_error),                   //         .error
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_0_reset_n),               // reset_in0.reset
		.clk            (clk_50_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_0_reset_n),                       // reset_in0.reset
		.clk            (sram_clk_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
